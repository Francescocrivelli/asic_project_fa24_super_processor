module ForwardingLogic(
    input [31:0] X_inst;
    input [31:0] D_inst;
    input [31:0] Mem_WB_inst;


);

always @(*) begin
    
end



endmodule
`include "const.vh"

module Riscv151(
    input clk,
    input reset,

    // Memory system ports
    output [31:0] dcache_addr,
    output [31:0] icache_addr,
    output [3:0] dcache_we,
    output dcache_re,
    output icache_re,
    output [31:0] dcache_din,
    input [31:0] dcache_dout,
    input [31:0] icache_dout,
    input stall,
    output [31:0] csr

);

  reg [31:0] PC;

  // Implement your core here, then delete this comment
  always @(*) begin
    if (reset) begin
      PC = PC_RESET;
      

    end
  end


endmodule
